// Osman Suzer
//
// 131044051
//

module _32_Bits_ALU_testbench();


	reg [31:0]a, b;
	reg [2:0] aluOp;
	
	wire c32;
	wire [31:0] r;
	wire Z, V;
	
	_32_Bits_ALU alu(r, c32, Z, V, a, b, aluOp);

	initial begin
	//and

	a =32'b00000000000000000000000000000000; 
	b =32'b00000000000000000000000000000000;
	aluOp = 3'b000;
	
	#10;
	a =32'b00000000000000000000000000000000; 
	b =32'b11111111111111111111111111111111;
	aluOp = 3'b000;
	
	#10;
	a =32'b11111111111111111111111111111111;
	b =32'b11111111111111111111111111111111;
	aluOp = 3'b000;
	
	//or
	#10;
	a =32'b00000000000000000000000000000000; 
	b =32'b00000000000000000000000000000000;
	aluOp = 3'b001;
	
	#10;
	a =32'b00000000000000000000000000000000; 
	b =32'b11111111111111111111111111111111;
	aluOp = 3'b001;
	
	#10;
	a =32'b11111111111111111111111111111111;
	b =32'b11111111111111111111111111111111;
	aluOp = 3'b001;
	
	
	// add
	
	#10;
	a =32'b00000000000000000000000000000000; 
	b =32'b00000000000000000000000000000000;
	aluOp = 3'b010;
	
	#10;
	a =32'b00000000000000000000000000000000; 
	b =32'b11111111111111111111111111111111;
	aluOp = 3'b010;
	
	#10;
	a =32'b11111111111111111111111111111111;
	b =32'b11111111111111111111111111111111;
	aluOp = 3'b010;
	

	//substract
	#10;
	a =32'b00000000000000000000000000000000; 
	b =32'b00000000000000000000000000000000;
	aluOp = 3'b110;
	
	#10;
	a =32'b00000000000000000000000000000000; 
	b =32'b01111111111111111111111111111111;
	aluOp = 3'b110;
	
	#10;
	a =32'b10000000000000000000000000000000; 
	b =32'b01111111111111111111111111111111;
	aluOp = 3'b110;
	
	#10;
	a =32'b11111111111111111111111111111111;
	b =32'b11111111111111111111111111111111;
	aluOp = 3'b110;
	
	#10;
	a =32'b00000000000000000000000000000100; 
	b =32'b00000000000000000000000000001010;
	aluOp = 3'b110;
	
	
	//set less than
	#10;
	a =32'b00000000000000000000000000000000; 
	b =32'b00000000000000000000000000000000;
	aluOp = 3'b111;
	
	#10;
	a =32'b00000000000000000000000000011000; 
	b =32'b00000000000000000000000000001111;
	aluOp = 3'b111;
	
	#10;
	a =32'b00000000000000000000000000000011; 
	b =32'b00000000000000000000000000001000;
	aluOp = 3'b111;
	
	#10;
	a =32'b00000000000000000000000000000000; 
	b =32'b11111111111111111111111111111111;
	aluOp = 3'b111;
	
	#10;
	a =32'b11111111111111111111111111111111;
	b =32'b11111111111111111111111111111111;
	aluOp = 3'b111;
	
	end
	
	initial begin
	$monitor("aluOp =>%3b a=%32b, b=%32b, result=%32b, c32=%1b, V=%1b, Z=%1b" , aluOp, a, b, r, c32, V, Z);
	end
	
	
endmodule